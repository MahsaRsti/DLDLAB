library verilog;
use verilog.vl_types.all;
entity wave_gen_core_tb is
end wave_gen_core_tb;
